module simula();

endmodule
