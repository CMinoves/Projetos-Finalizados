module ula (ALUctl, A, B,ALUOut, Zero);
input [3:0]ALUctl;
input [7:0] A,B;
output reg[7:0]ALUOut;
output Zero;
always @(ALUctl, A, B, Zero) begin //reevaluate if these change
case (ALUctl)
	1:ALUOut <= A/2;//hlf
	2:ALUOut <=A;//lfh
	3:Zero<= A == B ? 0 : 1; //bne
	4:ALUOut<= A//lw
	5:ALUOut<= A//sw
	6:Zero<= A == B ? 1 : 0; //beq
	7:ALUOut <= A+B; //cnt
	8:ALUOut <=B //set

default:ALUOut<= 0;
endcase
end
endmodule