library verilog;
use verilog.vl_types.all;
entity Contador3bits is
    port(
        clock           : in     vl_logic;
        reset           : in     vl_logic;
        num             : out    vl_logic_vector(2 downto 0)
    );
end Contador3bits;
