module processador(clock, operacao, tag, saidabus);
/*input clock;
input [1:0] operacao;
input [2:0] tag;
reg [9:0] b0,b1,b2,b3;
/*
	9-8: estado
	7-5: tag
	4-0: valor
*/


	
endmodule
