library verilog;
use verilog.vl_types.all;
entity decodificadorMARAvilhoso is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        l1              : out    vl_logic;
        l2              : out    vl_logic;
        l3              : out    vl_logic;
        l4              : out    vl_logic;
        l5              : out    vl_logic;
        l6              : out    vl_logic;
        l7              : out    vl_logic
    );
end decodificadorMARAvilhoso;
