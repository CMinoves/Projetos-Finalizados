library verilog;
use verilog.vl_types.all;
entity processor is
    port(
        DIN             : in     vl_logic_vector(15 downto 0);
        Resetn          : in     vl_logic;
        Clock           : in     vl_logic;
        Run             : in     vl_logic;
        Done            : out    vl_logic;
        \Bus\           : out    vl_logic_vector(15 downto 0)
    );
end processor;
